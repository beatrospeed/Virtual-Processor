library verilog;
use verilog.vl_types.all;
entity div_testbench is
end div_testbench;
