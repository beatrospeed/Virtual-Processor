library verilog;
use verilog.vl_types.all;
entity SelectEncode is
    port(
        R0in            : out    vl_logic_vector(15 downto 0);
        R1in            : out    vl_logic_vector(15 downto 0);
        R2in            : out    vl_logic_vector(15 downto 0);
        R3in            : out    vl_logic_vector(15 downto 0);
        R4in            : out    vl_logic_vector(15 downto 0);
        R5in            : out    vl_logic_vector(15 downto 0);
        R6in            : out    vl_logic_vector(15 downto 0);
        R7in            : out    vl_logic_vector(15 downto 0);
        R8in            : out    vl_logic_vector(15 downto 0);
        R9in            : out    vl_logic_vector(15 downto 0);
        R10in           : out    vl_logic_vector(15 downto 0);
        R11in           : out    vl_logic_vector(15 downto 0);
        R12in           : out    vl_logic_vector(15 downto 0);
        R13in           : out    vl_logic_vector(15 downto 0);
        R14in           : out    vl_logic_vector(15 downto 0);
        R15in           : out    vl_logic_vector(15 downto 0);
        R0out           : out    vl_logic_vector(15 downto 0);
        R1out           : out    vl_logic_vector(15 downto 0);
        R2out           : out    vl_logic_vector(15 downto 0);
        R3out           : out    vl_logic_vector(15 downto 0);
        R4out           : out    vl_logic_vector(15 downto 0);
        R5out           : out    vl_logic_vector(15 downto 0);
        R6out           : out    vl_logic_vector(15 downto 0);
        R7out           : out    vl_logic_vector(15 downto 0);
        R8out           : out    vl_logic_vector(15 downto 0);
        R9out           : out    vl_logic_vector(15 downto 0);
        R10out          : out    vl_logic_vector(15 downto 0);
        R11out          : out    vl_logic_vector(15 downto 0);
        R12out          : out    vl_logic_vector(15 downto 0);
        R13out          : out    vl_logic_vector(15 downto 0);
        R14out          : out    vl_logic_vector(15 downto 0);
        R15out          : out    vl_logic_vector(15 downto 0);
        c_sign_extended : out    vl_logic_vector(31 downto 0);
        IRin            : in     vl_logic_vector(31 downto 0);
        Rin             : in     vl_logic;
        Rout            : in     vl_logic;
        BAout           : in     vl_logic;
        GRA             : in     vl_logic;
        GRB             : in     vl_logic;
        GRC             : in     vl_logic
    );
end SelectEncode;
