library verilog;
use verilog.vl_types.all;
entity dataPath is
    port(
        PCout           : in     vl_logic;
        Zlowout         : in     vl_logic;
        MDRout          : in     vl_logic;
        R2out           : in     vl_logic;
        R4out           : in     vl_logic;
        MARin           : in     vl_logic;
        Zin             : in     vl_logic;
        PCin            : in     vl_logic;
        MDRin           : in     vl_logic;
        IRin            : in     vl_logic;
        Yin             : in     vl_logic;
        IncPc           : in     vl_logic;
        read            : in     vl_logic;
        R5in            : in     vl_logic;
        R2in            : in     vl_logic;
        R4in            : in     vl_logic;
        clk             : in     vl_logic;
        control         : in     vl_logic_vector(3 downto 0);
        Mdatain         : in     vl_logic_vector(31 downto 0);
        R0out           : in     vl_logic;
        R1out           : in     vl_logic;
        R3out           : in     vl_logic;
        R5out           : in     vl_logic;
        R6out           : in     vl_logic;
        R7out           : in     vl_logic;
        R8out           : in     vl_logic;
        R9out           : in     vl_logic;
        R10out          : in     vl_logic;
        R11out          : in     vl_logic;
        R12out          : in     vl_logic;
        R13out          : in     vl_logic;
        R14out          : in     vl_logic;
        R15out          : in     vl_logic;
        HIout           : in     vl_logic;
        LOout           : in     vl_logic;
        InPortout       : in     vl_logic;
        OutPortout      : in     vl_logic;
        Cout            : in     vl_logic;
        Zhighout        : in     vl_logic;
        R0in            : in     vl_logic;
        R1in            : in     vl_logic;
        R3in            : in     vl_logic;
        R6in            : in     vl_logic;
        R7in            : in     vl_logic;
        R8in            : in     vl_logic;
        R9in            : in     vl_logic;
        R10in           : in     vl_logic;
        R11in           : in     vl_logic;
        R12in           : in     vl_logic;
        R13in           : in     vl_logic;
        R14in           : in     vl_logic;
        R15in           : in     vl_logic;
        HIin            : in     vl_logic;
        LOin            : in     vl_logic;
        Zhighin         : in     vl_logic;
        Zlowin          : in     vl_logic;
        InPortin        : in     vl_logic;
        Cin             : in     vl_logic;
        reset           : in     vl_logic;
        R0Val           : out    vl_logic_vector(31 downto 0);
        R1Val           : out    vl_logic_vector(31 downto 0);
        R2Val           : out    vl_logic_vector(31 downto 0);
        R3Val           : out    vl_logic_vector(31 downto 0);
        R4Val           : out    vl_logic_vector(31 downto 0);
        R5Val           : out    vl_logic_vector(31 downto 0);
        R6Val           : out    vl_logic_vector(31 downto 0);
        R7Val           : out    vl_logic_vector(31 downto 0);
        R8Val           : out    vl_logic_vector(31 downto 0);
        R9Val           : out    vl_logic_vector(31 downto 0);
        R10Val          : out    vl_logic_vector(31 downto 0);
        R11Val          : out    vl_logic_vector(31 downto 0);
        R12Val          : out    vl_logic_vector(31 downto 0);
        R13Val          : out    vl_logic_vector(31 downto 0);
        R14Val          : out    vl_logic_vector(31 downto 0);
        R15Val          : out    vl_logic_vector(31 downto 0);
        \bus\           : out    vl_logic_vector(31 downto 0)
    );
end dataPath;
