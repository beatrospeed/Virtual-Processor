library verilog;
use verilog.vl_types.all;
entity dataPath is
    port(
        PCout           : in     vl_logic;
        Zlowout         : in     vl_logic;
        MDRout          : in     vl_logic;
        MARin           : in     vl_logic;
        Zin             : in     vl_logic;
        PCin            : in     vl_logic;
        MDRin           : in     vl_logic;
        read            : in     vl_logic;
        write           : in     vl_logic;
        IRin            : in     vl_logic;
        Yin             : in     vl_logic;
        IncPc           : in     vl_logic;
        clk             : in     vl_logic;
        mdr_read        : in     vl_logic_vector(1 downto 0);
        control         : in     vl_logic_vector(3 downto 0);
        HIout           : in     vl_logic;
        LOout           : in     vl_logic;
        InPortout       : in     vl_logic;
        OutPortout      : in     vl_logic;
        Cout            : in     vl_logic;
        Zhighout        : in     vl_logic;
        HIin            : in     vl_logic;
        LOin            : in     vl_logic;
        Zhighin         : in     vl_logic;
        Zlowin          : in     vl_logic;
        InPortin        : in     vl_logic;
        Cin             : in     vl_logic;
        reset           : in     vl_logic;
        BAout           : in     vl_logic;
        OutPortin       : in     vl_logic;
        Rin             : in     vl_logic;
        Rout            : in     vl_logic;
        GRA             : in     vl_logic;
        GRB             : in     vl_logic;
        GRC             : in     vl_logic;
        Immediate       : in     vl_logic_vector(31 downto 0);
        R0Val           : out    vl_logic_vector(31 downto 0);
        R1Val           : out    vl_logic_vector(31 downto 0);
        R2Val           : out    vl_logic_vector(31 downto 0);
        R3Val           : out    vl_logic_vector(31 downto 0);
        R4Val           : out    vl_logic_vector(31 downto 0);
        R5Val           : out    vl_logic_vector(31 downto 0);
        R6Val           : out    vl_logic_vector(31 downto 0);
        R7Val           : out    vl_logic_vector(31 downto 0);
        R8Val           : out    vl_logic_vector(31 downto 0);
        R9Val           : out    vl_logic_vector(31 downto 0);
        R10Val          : out    vl_logic_vector(31 downto 0);
        R11Val          : out    vl_logic_vector(31 downto 0);
        R12Val          : out    vl_logic_vector(31 downto 0);
        R13Val          : out    vl_logic_vector(31 downto 0);
        R14Val          : out    vl_logic_vector(31 downto 0);
        R15Val          : out    vl_logic_vector(31 downto 0);
        IRval           : out    vl_logic_vector(31 downto 0);
        \bus\           : out    vl_logic_vector(31 downto 0);
        MDRval          : out    vl_logic_vector(31 downto 0);
        mux_data_out    : out    vl_logic_vector(31 downto 0);
        YVal            : out    vl_logic_vector(31 downto 0);
        R0TempOut       : out    vl_logic_vector(31 downto 0);
        C_sign_extended : out    vl_logic_vector(31 downto 0);
        InPort_D        : out    vl_logic_vector(31 downto 0);
        OutPort_D       : out    vl_logic_vector(31 downto 0);
        PCVal           : out    vl_logic_vector(31 downto 0);
        CVal            : out    vl_logic_vector(31 downto 0);
        Mdatain         : out    vl_logic_vector(31 downto 0);
        ZVal            : out    vl_logic_vector(63 downto 0);
        ALUVal_D        : out    vl_logic_vector(63 downto 0);
        Rin_Select      : out    vl_logic_vector(15 downto 0);
        Rout_Select     : out    vl_logic_vector(15 downto 0);
        MAR_D           : out    vl_logic_vector(31 downto 0)
    );
end dataPath;
