library verilog;
use verilog.vl_types.all;
entity dataPath is
    port(
        R0in            : in     vl_logic;
        R1in            : in     vl_logic;
        R2in            : in     vl_logic;
        R3in            : in     vl_logic;
        R4in            : in     vl_logic;
        R5in            : in     vl_logic;
        R6in            : in     vl_logic;
        R7in            : in     vl_logic;
        R8in            : in     vl_logic;
        R9in            : in     vl_logic;
        R10in           : in     vl_logic;
        R11in           : in     vl_logic;
        R12in           : in     vl_logic;
        R13in           : in     vl_logic;
        R14in           : in     vl_logic;
        R15in           : in     vl_logic;
        Yin             : in     vl_logic;
        Zin             : in     vl_logic;
        HIin            : in     vl_logic;
        LOin            : in     vl_logic;
        InPortin        : in     vl_logic;
        OutPortin       : in     vl_logic;
        MARin           : in     vl_logic;
        MDRin           : in     vl_logic;
        IRin            : in     vl_logic;
        PCin            : in     vl_logic;
        BusMuxin_R0     : out    vl_logic;
        BusMuxin_R1     : out    vl_logic;
        BusMuxin_R2     : out    vl_logic;
        BusMuxin_R3     : out    vl_logic;
        BusMuxin_R4     : out    vl_logic;
        BusMuxin_R5     : out    vl_logic;
        BusMuxin_R6     : out    vl_logic;
        BusMuxin_R7     : out    vl_logic;
        BusMuxin_R8     : out    vl_logic;
        BusMuxin_R9     : out    vl_logic;
        BusMuxin_R10    : out    vl_logic;
        BusMuxin_R11    : out    vl_logic;
        BusMuxin_R12    : out    vl_logic;
        BusMuxin_R13    : out    vl_logic;
        BusMuxin_R14    : out    vl_logic;
        BusMuxin_R15    : out    vl_logic;
        BusMuxin_HIout  : out    vl_logic;
        BusMuxin_LOout  : out    vl_logic;
        BusMuxin_Zhighout: out    vl_logic;
        BusMuxin_Zlowout: out    vl_logic;
        BusMuxin_PCout  : out    vl_logic;
        BusMuxin_MDRout : out    vl_logic;
        BusMuxin_In_Portout: out    vl_logic;
        BusMuxin_Cin    : out    vl_logic;
        BusMuxin_in24   : out    vl_logic;
        BusMuxin_in25   : out    vl_logic;
        BusMuxin_in26   : out    vl_logic;
        BusMuxin_in27   : out    vl_logic;
        BusMuxin_in28   : out    vl_logic;
        BusMuxin_in29   : out    vl_logic;
        BusMuxin_in30   : out    vl_logic;
        BusMuxin_in31   : out    vl_logic;
        Y_in            : out    vl_logic;
        Z_in            : out    vl_logic;
        R0Val           : out    vl_logic_vector(31 downto 0);
        R1Val           : out    vl_logic_vector(31 downto 0);
        R2Val           : out    vl_logic_vector(31 downto 0);
        R3Val           : out    vl_logic_vector(31 downto 0);
        R4Val           : out    vl_logic_vector(31 downto 0);
        R5Val           : out    vl_logic_vector(31 downto 0);
        R6Val           : out    vl_logic_vector(31 downto 0);
        R7Val           : out    vl_logic_vector(31 downto 0);
        R8Val           : out    vl_logic_vector(31 downto 0);
        R9Val           : out    vl_logic_vector(31 downto 0);
        R10Val          : out    vl_logic_vector(31 downto 0);
        R11Val          : out    vl_logic_vector(31 downto 0);
        R12Val          : out    vl_logic_vector(31 downto 0);
        R13Val          : out    vl_logic_vector(31 downto 0);
        R14Val          : out    vl_logic_vector(31 downto 0);
        R15Val          : out    vl_logic_vector(31 downto 0);
        load            : in     vl_logic;
        clk             : in     vl_logic;
        reset           : in     vl_logic;
        Mdata_in        : in     vl_logic_vector(31 downto 0);
        control         : in     vl_logic_vector(3 downto 0);
        ADD             : in     vl_logic;
        SUB             : in     vl_logic;
        MUL             : in     vl_logic;
        DIV             : in     vl_logic;
        SHR             : in     vl_logic;
        SHL             : in     vl_logic;
        \ROR\           : in     vl_logic;
        \ROL\           : in     vl_logic;
        \AND\           : in     vl_logic;
        \OR\            : in     vl_logic;
        NEG             : in     vl_logic;
        \NOT\           : in     vl_logic;
        IncPc           : in     vl_logic;
        Mdatain         : out    vl_logic_vector(31 downto 0);
        ZVal            : out    vl_logic_vector(63 downto 0);
        \bus\           : out    vl_logic_vector(31 downto 0);
        IRval           : out    vl_logic_vector(31 downto 0);
        MDRval          : out    vl_logic_vector(31 downto 0);
        HIval           : out    vl_logic_vector(31 downto 0);
        LOval           : out    vl_logic_vector(31 downto 0)
    );
end dataPath;
