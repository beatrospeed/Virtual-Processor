module RAM (output reg [31:0] RAMout/* to MDR MDataIN*/, input read, input write,input [31:0] data/*FROm MDR AKA Q*/, input [8:0] Address/*From MAR*/);



endmodule