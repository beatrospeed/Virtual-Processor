library verilog;
use verilog.vl_types.all;
entity Mux_32_to_1 is
    port(
        BusMuxOut       : out    vl_logic_vector(31 downto 0);
        \Select\        : in     vl_logic_vector(4 downto 0);
        BusMuxin_R0     : in     vl_logic;
        BusMuxin_R1     : in     vl_logic;
        BusMuxin_R2     : in     vl_logic;
        BusMuxin_R3     : in     vl_logic;
        BusMuxin_R4     : in     vl_logic;
        BusMuxin_R5     : in     vl_logic;
        BusMuxin_R6     : in     vl_logic;
        BusMuxin_R7     : in     vl_logic;
        BusMuxin_R8     : in     vl_logic;
        BusMuxin_R9     : in     vl_logic;
        BusMuxin_R10    : in     vl_logic;
        BusMuxin_R11    : in     vl_logic;
        BusMuxin_R12    : in     vl_logic;
        BusMuxin_R13    : in     vl_logic;
        BusMuxin_R14    : in     vl_logic;
        BusMuxin_R15    : in     vl_logic;
        BusMuxin_HIout  : in     vl_logic;
        BusMuxin_LOout  : in     vl_logic;
        BusMuxin_Zhighout: in     vl_logic;
        BusMuxin_Zlowout: in     vl_logic;
        BusMuxin_PCout  : in     vl_logic;
        BusMuxin_MDRout : in     vl_logic;
        BusMuxin_In_Portout: in     vl_logic;
        BusMuxin_Cout   : in     vl_logic;
        BusMuxin_in24   : in     vl_logic;
        BusMuxin_in25   : in     vl_logic;
        BusMuxin_in26   : in     vl_logic;
        BusMuxin_in27   : in     vl_logic;
        BusMuxin_in28   : in     vl_logic;
        BusMuxin_in29   : in     vl_logic;
        BusMuxin_in30   : in     vl_logic;
        BusMuxin_in31   : in     vl_logic
    );
end Mux_32_to_1;
